library verilog;
use verilog.vl_types.all;
entity edt_top_blockB_v_ctl is
end edt_top_blockB_v_ctl;
