library verilog;
use verilog.vl_types.all;
entity dff_sr_0 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end dff_sr_0;
