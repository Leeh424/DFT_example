library verilog;
use verilog.vl_types.all;
entity latch_s is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end latch_s;
