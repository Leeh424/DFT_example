library verilog;
use verilog.vl_types.all;
entity inv16 is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end inv16;
