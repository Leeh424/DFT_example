library verilog;
use verilog.vl_types.all;
entity trib08 is
    port(
        A               : in     vl_logic;
        E               : in     vl_logic;
        Y               : out    vl_logic
    );
end trib08;
