library verilog;
use verilog.vl_types.all;
entity buf02 is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end buf02;
