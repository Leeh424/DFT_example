library verilog;
use verilog.vl_types.all;
entity and02 is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        Y               : out    vl_logic
    );
end and02;
