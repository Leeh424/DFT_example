library verilog;
use verilog.vl_types.all;
entity aoi332 is
    port(
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        Y               : out    vl_logic
    );
end aoi332;
